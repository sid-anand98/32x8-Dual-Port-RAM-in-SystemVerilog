parameter ADDR_WIDTH=4;
parameter DATA_WIDTH=7;
parameter MEM_SIZE=31;
